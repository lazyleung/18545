module interrupt(
        clock, reset,
        IF_in, IE_in, IF_load, IE_load
    );


endmodule // interrupt