module oamram_test(
		   I_MEM_CLK,
		   I_RESET,
		   I_OAM_ADDR,
		   IO_OAM_DATA,
		   I_OAM_WE_L,
		   I_OAM_RE_L
		   );

   input        I_MEM_CLK, I_RESET;
   input [15:0] I_OAM_ADDR;
   inout [7:0] 	IO_OAM_DATA;
   input 	    I_OAM_WE_L, I_OAM_RE_L;
   
   wire 	bram_en;
   wire 	bram_we;
   wire [15:0] 	router_addr;
   wire [15:0] 	bram_banked_addr;
   wire [15:0] 	bram_addr;
   wire [7:0] 	bram_data_in2, bram_data_out2;
   
   assign bram_addr = router_addr[14:0];
   

   bram_wrapper #(16'h00FF) ifconverter(
				       .I_CLK(I_MEM_CLK),
				       .I_RESET(I_RESET),
				       .I_ADDR(I_OAM_ADDR),
				       .IO_DATA(IO_OAM_DATA),
				       .I_WE_L(I_OAM_WE_L),
				       .I_RE_L(I_OAM_RE_L),
				       .O_BRAM_EN(bram_en),
				       .O_BRAM_WE(bram_we),
				       .O_BRAM_ADDR(router_addr),
				       .O_BRAM_DIN(bram_data_in2),
				       .I_BRAM_DOUT(bram_data_out2)
				       );


      /* Actual Memory Location*/
   bram_lcd lcdbram(
		.clka(I_MEM_CLK),
		.wea(bram_we),
		.addra(bram_addr),
		.dina(bram_data_in2),
		.douta(bram_data_out2)
		);

   
endmodule 