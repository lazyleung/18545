module interrupt(
        I_CLOCK, I_RESET,
        IF_in, IE_in, IF_load, IE_load
    );


endmodule // interrupt