module squarewave_generator(
                            /*System Level Inputs*/
                            I_BITCLK,
                            I_RESET,

			    /*Sampling Strobe Input*/
			    I_STROBE,
			    
                            /*Waveform Output Signal*/
                            O_SAMPLE,
			    
                            /*User Freq & Duty Cycle Spec*/
                            I_FREQUENCY,
                            I_DUTY_CYCLE,
                            I_WAVEFORM_EN, 
			    I_VOLUME);
   
   
   input I_BITCLK, I_RESET;
   output reg [19:0] O_SAMPLE;
   input 	     I_WAVEFORM_EN, I_STROBE;
   input [10:0]      I_FREQUENCY; //will be calculated as 2^17/(2^11-I_FREQUENCY)
   input [3:0] 	     I_VOLUME;
   input [1:0] 	     I_DUTY_CYCLE; /* 00 - 12.5%
				    * 01 - 25%
				    * 10 - 50%
				    * 11 - 75% */
   
   wire [15:0] 	     num_strobes_in_period;
   wire [15:0] 	     num_strobes_high;
   reg [10:0] 	     freq_reg, freq_reg_d1, freq_reg_d2;
   reg [1:0] 	     duty_cyc_reg, duty_cyc_reg_d1, duty_cyc_reg_d2;
   reg [3:0] 	     volume_reg, volume_reg_d1, volume_reg_d2;
   reg 		     waveform;
   reg [15:0] 	     count;

   wire [19:0] 	     volume_to_sample;
   
   /*go from a 4 bit value to a 20 bit value*/
   assign volume_to_sample = volume_reg << 16;
   
   /*figure out the duty cycle*/
   assign num_strobes_high = (duty_cyc_reg == 'b00) ? num_strobes_in_period >> 3 : //12.5%
                             (duty_cyc_reg == 'b01) ? num_strobes_in_period >> 2 : //25%
                             (duty_cyc_reg == 'b10) ? num_strobes_in_period >> 1 : //50%
                             (duty_cyc_reg == 'b11) ? (num_strobes_in_period + //75%
						       num_strobes_in_period << 1) >> 2 
			     : 0; 

   /* Cross information over clock domains by
    * registering the information a few times*/
   always @(posedge I_BITCLK) begin
      freq_reg_d1 <= I_FREQUENCY;
      duty_cyc_reg_d1 <= I_DUTY_CYCLE;
      volume_reg_d1 <= I_VOLUME;
      freq_reg_d2 <= freq_reg_d1;
      duty_cyc_reg_d2 <= duty_cyc_reg_d1;
      volume_reg_d2 <= volume_reg_d1;
      freq_reg <= freq_reg_d2;
      duty_cyc_reg <= duty_cyc_reg_d2;
      volume_reg <= volume_reg_d2;
   end

   /*generate the square waveform based on the specification*/
   always @(posedge I_BITCLK) begin

      if (I_STROBE) begin
			count <= count + 1;
	 
			/*make the duty cycle*/
			//if (count < num_strobes_high) begin
			if (count < 48000/880) begin
            O_SAMPLE <= 20'h80000;
			end
	 
			/*low end of duty cycle, finish period*/
			//else if (count < num_strobes_in_period) begin
			else if (count < 48000/440) begin
            O_SAMPLE <= 20'h7ffff;
			end
	 
			/*reset the counter when overflow*/
			//else if (count >= num_strobes_in_period) begin
			else if (count >= 48000/440) begin
            count <= 0;
			end
	 
		end // if (I_STROBE)

      /*If not enabled, disable the output*/
      //if (~I_WAVEFORM_EN)
			//O_SAMPLE <= 0;

      if (I_RESET) begin
         count <= 0;
			O_SAMPLE <= 0;
      end
      
   end // always @ (posedge I_BITCLK)
      
   wire gnd = 0;

   /* Translate the frequency to the strobes in period
    * from the BRAM lookup table*/
   sound_bram period_lookup_table(
		                  .clka(I_BITCLK),
		                  .wea(gnd),
		                  .addra(freq_reg),
		                  .dina(0),
		                  .douta(num_strobes_in_period)
		                  );
   


endmodule