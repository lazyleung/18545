`define CARTRIDGE_LO 'h0000
`define CARTRIDGE_HI 'h7fff

`define EXTERNAL_EXPANSION_LO 'hA000
`define EXTERNAL_EXPANSION_HI 'hBFFF

`define LCDRAM_LO 'h8000
`define LCDRAM_HI 'h9FFF

`define WRAM_LO 'hC000
`define WRAM_HI 'hCFFF

`define OAM_LO 'hFE00
`define OAM_HI 'hFF7F

`define LWRAM_LO 'hFF80
`define LWRAM_HI 'hFFFE

`define IOREG_LO 'hFF00
`define IOREG_HI 'hFF7F

`define IE_REGISTER 'hFFFF